module Random_Circuit_7 (
    input A, B, clk, rst,
    output reg Q
);
    wire or_out, nand_out, xor_out;
    
    or (or_out, A, B);
    nand (nand_out, A, B);
    xor (xor_out, A, B);
    
    always @(posedge clk or posedge rst) begin
        if (rst)
            Q <= 0;
        else
            Q <= or_out | nand_out ^ xor_out;
    end
endmodule
