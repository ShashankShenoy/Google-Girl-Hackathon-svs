module nand_buffer_flipflop (
    input wire clk,
    input wire rst,
    input wire a,
    input wire b,
    output reg q
);

wire nand_out, buf_out;

assign nand_out = ~(a & b); // NAND gate
assign buf_out = nand_out;  // Buffer

always @(posedge clk or posedge rst) begin
    if (rst)
        q <= 0;
    else
        q <= buf_out;
end

endmodule
